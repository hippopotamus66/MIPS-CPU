    Mac OS X            	   2   �                                           ATTR         �   L                  �     com.apple.lastuseddate#PS       �   <  com.apple.quarantine O��]    ww�    q/0081;5fa20612;Chrome;6646E9C7-4D1B-4F56-9206-E6B366C022D1 