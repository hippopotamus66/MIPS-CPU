library ieee;
use ieee.std_logic_1164.all;
use work.eecs361_gates.all;
use ieee.numeric_std.all; 
use ieee.std_logic_arith.all;
use work.eecs361.mux_n;
use ieee.std_logic_signed.all;
entity sll_32bit is
port (
  	x     : in std_logic_vector(31 downto 0);
   	shift     : in std_logic_vector(31 downto 0);
   	--cin   : in std_logic;
     	z     : out std_logic_vector(31 downto 0)
    	--cout  : out std_logic
);
end sll_32bit;
architecture structural of sll_32bit is
signal xin : std_logic_vector(31 downto 0);
signal test : std_logic_vector(0 to 31);
signal t : std_logic_vector(31 downto 0);
	component mux_32to1 is
		  port (
			sel   : in  std_logic_vector(4 downto 0);
			src  : in  std_logic_vector(31 downto 0);
			z	    : out std_logic
  			);
        end component;
begin
xin <= "00000000000000000000000000000000";
test (0 to 31) <= x(31 downto 0);
 	 mux_map0: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(0),
				src(31 downto 1) => xin(31 downto 1),
	  			z => z(0)
				);
 	 mux_map1: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(1),
				src(1) => x(0),
				src(31 downto 2) => xin(31 downto 2),
	  			z => z(1)
				);
 	 mux_map2: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(2),
				src(1) => x(1),
				src(2) => x(0),
				src(31 downto 3) => xin(31 downto 3),
	  			z => z(2)
				);
 	 mux_map3: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(3),
				src(1) => x(2),
				src(2) => x(1),
				src(3) => x(0),
				src(31 downto 4) => xin(31 downto 4),
	  			z => z(3)
				);
 	 mux_map4: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(4),
				src(1) => x(3),
				src(2) => x(2),
				src(3) => x(1),
				src(4) => x(0),
				src(31 downto 5) => xin(31 downto 5),
	  			z => z(4)
				);
 	 mux_map5: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(5),
				src(1) => x(4),
				src(2) => x(3),
				src(3) => x(3),
				src(4) => x(1),
				src(5) => x(0),
				src(31 downto 6) => xin(31 downto 6),
	  			z => z(5)
				);
 	 mux_map6: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(6),
				src(1) => x(5),
				src(2) => x(4),
				src(3) => x(3),
				src(4) => x(2),
				src(5) => x(1),
				src(6) => x(0),
				src(31 downto 7) => xin(31 downto 7),
	  			z => z(6)
				);
 	 mux_map7: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(7),
				src(1) => x(6),
				src(2) => x(5),
				src(3) => x(4),
				src(4) => x(3),
				src(5) => x(2),
				src(6) => x(1),
				src(7) => x(0),
				src(31 downto 8) => xin(31 downto 8),
	  			z => z(7)
				);
 	 mux_map8: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(8),
				src(1) => x(7),
				src(2) => x(6),
				src(3) => x(5),
				src(4) => x(4),
				src(5) => x(3),
				src(6) => x(2),
				src(7) => x(1),
				src(8) => x(0),
				src(31 downto 9) => xin(31 downto 9),
	  			z => z(8)
				);
 	 mux_map9: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(9),
				src(1) => x(8),
				src(2) => x(7),
				src(3) => x(6),
				src(4) => x(5),
				src(5) => x(4),
				src(6) => x(3),
				src(7) => x(2),
				src(8) => x(1),
				src(9) => x(0),
				src(31 downto 10) => xin(31 downto 10),
	  			z => z(9)
				);
 	 mux_map10: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(10),
				src(1) => x(9),
				src(2) => x(8),
				src(3) => x(7),
				src(4) => x(6),
				src(5) => x(5),
				src(6) => x(4),
				src(7) => x(3),
				src(8) => x(2),
				src(9) => x(1),
				src(10) => x(0),
				src(31 downto 11) => xin(31 downto 11),
	  			z => z(10)
				);
 	 mux_map11: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(11),
				src(1) => x(10),
				src(2) => x(9),
				src(3) => x(8),
				src(4) => x(7),
				src(5) => x(6),
				src(6) => x(5),
				src(7) => x(4),
				src(8) => x(3),
				src(9) => x(2),
				src(10) => x(1),
				src(11) => x(0),
				src(31 downto 12) => xin(31 downto 12),
	  			z => z(11)
				);
 	 mux_map12: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(12),
				src(1) => x(11),
				src(2) => x(10),
				src(3) => x(9),
				src(4) => x(8),
				src(5) => x(7),
				src(6) => x(6),
				src(7) => x(5),
				src(8) => x(4),
				src(9) => x(3),
				src(10) => x(2),
				src(11) => x(1),
				src(12) => x(0),
				src(31 downto 13) => xin(31 downto 13),
	  			z => z(12)
				);
 	 mux_map13: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(13),
				src(1) => x(12),
				src(2) => x(11),
				src(3) => x(10),
				src(4) => x(9),
				src(5) => x(8),
				src(6) => x(7),
				src(7) => x(6),
				src(8) => x(5),
				src(9) => x(4),
				src(10) => x(3),
				src(11) => x(2),
				src(12) => x(1),
				src(13) => x(0),
				src(31 downto 14) => xin(31 downto 14),
	  			z => z(13)
				);
 	 mux_map14: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(14),
				src(1) => x(13),
				src(2) => x(12),
				src(3) => x(11),
				src(4) => x(10),
				src(5) => x(9),
				src(6) => x(8),
				src(7) => x(7),
				src(8) => x(6),
				src(9) => x(5),
				src(10) => x(4),
				src(11) => x(3),
				src(12) => x(2),
				src(13) => x(1),
				src(14) => x(0),
				src(31 downto 15) => xin(31 downto 15),
	  			z => z(14)
				);
 	 mux_map15: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(15),
				src(1) => x(14),
				src(2) => x(13),
				src(3) => x(12),
				src(4) => x(11),
				src(5) => x(10),
				src(6) => x(9),
				src(7) => x(8),
				src(8) => x(7),
				src(9) => x(6),
				src(10) => x(5),
				src(11) => x(4),
				src(12) => x(3),
				src(13) => x(2),
				src(14) => x(1),
				src(15) => x(0),
				src(31 downto 16) => xin(31 downto 16),
	  			z => z(15)
				);
 	 mux_map16: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(16),
				src(1) => x(15),
				src(2) => x(14),
				src(3) => x(13),
				src(4) => x(12),
				src(5) => x(11),
				src(6) => x(10),
				src(7) => x(9),
				src(8) => x(8),
				src(9) => x(7),
				src(10) => x(6),
				src(11) => x(5),
				src(12) => x(4),
				src(13) => x(3),
				src(14) => x(2),
				src(15) => x(1),
				src(16) => x(0),
				src(31 downto 17) => xin(31 downto 17),
	  			z => z(16)
				);
 	 mux_map17: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(17),
				src(1) => x(16),
				src(2) => x(15),
				src(3) => x(14),
				src(4) => x(13),
				src(5) => x(12),
				src(6) => x(11),
				src(7) => x(10),
				src(8) => x(9),
				src(9) => x(8),
				src(10) => x(7),
				src(11) => x(6),
				src(12) => x(5),
				src(13) => x(4),
				src(14) => x(3),
				src(15) => x(2),
				src(16) => x(1),
				src(17) => x(0),
				src(31 downto 18) => xin(31 downto 18),
	  			z => z(17)
				);
 	 mux_map18: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(18),
				src(1) => x(17),
				src(2) => x(16),
				src(3) => x(15),
				src(4) => x(14),
				src(5) => x(13),
				src(6) => x(12),
				src(7) => x(11),
				src(8) => x(10),
				src(9) => x(9),
				src(10) => x(8),
				src(11) => x(7),
				src(12) => x(6),
				src(13) => x(5),
				src(14) => x(4),
				src(15) => x(3),
				src(16) => x(2),
				src(17) => x(1),
				src(18) => x(0),
				src(31 downto 19) => xin(31 downto 19),
	  			z => z(18)
				);
 	 mux_map19: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(19),
				src(1) => x(18),
				src(2) => x(17),
				src(3) => x(16),
				src(4) => x(15),
				src(5) => x(14),
				src(6) => x(13),
				src(7) => x(12),
				src(8) => x(11),
				src(9) => x(10),
				src(10) => x(9),
				src(11) => x(8),
				src(12) => x(7),
				src(13) => x(6),
				src(14) => x(5),
				src(15) => x(4),
				src(16) => x(3),
				src(17) => x(2),
				src(18) => x(1),
				src(19) => x(0),
				src(31 downto 20) => xin(31 downto 20),
	  			z => z(19)
				);
 	 mux_map20: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(20),
				src(1) => x(19),
				src(2) => x(18),
				src(3) => x(17),
				src(4) => x(16),
				src(5) => x(15),
				src(6) => x(14),
				src(7) => x(13),
				src(8) => x(12),
				src(9) => x(11),
				src(10) => x(10),
				src(11) => x(9),
				src(12) => x(8),
				src(13) => x(7),
				src(14) => x(6),
				src(15) => x(5),
				src(16) => x(4),
				src(17) => x(3),
				src(18) => x(2),
				src(19) => x(1),
				src(20) => x(0),
				src(31 downto 21) => xin(31 downto 21),
	  			z => z(20)
				);
 	 mux_map21: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(21),
				src(1) => x(20),
				src(2) => x(19),
				src(3) => x(18),
				src(4) => x(17),
				src(5) => x(16),
				src(6) => x(15),
				src(7) => x(14),
				src(8) => x(13),
				src(9) => x(12),
				src(10) => x(11),
				src(11) => x(10),
				src(12) => x(9),
				src(13) => x(8),
				src(14) => x(7),
				src(15) => x(6),
				src(16) => x(5),
				src(17) => x(4),
				src(18) => x(3),
				src(19) => x(2),
				src(20) => x(1),
				src(21) => x(0),
				src(31 downto 22) => xin(31 downto 22),
	  			z => z(21)
				);
 	mux_map22: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(22),
				src(1) => x(21),
				src(2) => x(20),
				src(3) => x(19),
				src(4) => x(18),
				src(5) => x(17),
				src(6) => x(16),
				src(7) => x(15),
				src(8) => x(14),
				src(9) => x(13),
				src(10) => x(12),
				src(11) => x(11),
				src(12) => x(10),
				src(13) => x(9),
				src(14) => x(8),
				src(15) => x(7),
				src(16) => x(6),
				src(17) => x(5),
				src(18) => x(4),
				src(19) => x(3),
				src(20) => x(2),
				src(21) => x(1),
				src(22) => x(0),
				src(31 downto 23) => xin(31 downto 23),
	  			z => z(22)
				);
 	mux_map23: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(23),
				src(1) => x(22),
				src(2) => x(21),
				src(3) => x(20),
				src(4) => x(19),
				src(5) => x(18),
				src(6) => x(17),
				src(7) => x(16),
				src(8) => x(15),
				src(9) => x(14),
				src(10) => x(13),
				src(11) => x(12),
				src(12) => x(11),
				src(13) => x(10),
				src(14) => x(9),
				src(15) => x(8),
				src(16) => x(7),
				src(17) => x(6),
				src(18) => x(5),
				src(19) => x(4),
				src(20) => x(3),
				src(21) => x(2),
				src(22) => x(1),
				src(23) => x(0),
				src(31 downto 24) => xin(31 downto 24),
	  			z => z(23)
				);
 	mux_map24: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(24),
				src(1) => x(23),
				src(2) => x(22),
				src(3) => x(21),
				src(4) => x(20),
				src(5) => x(19),
				src(6) => x(18),
				src(7) => x(17),
				src(8) => x(16),
				src(9) => x(15),
				src(10) => x(14),
				src(11) => x(13),
				src(12) => x(12),
				src(13) => x(11),
				src(14) => x(10),
				src(15) => x(9),
				src(16) => x(8),
				src(17) => x(7),
				src(18) => x(6),
				src(19) => x(5),
				src(20) => x(4),
				src(21) => x(3),
				src(22) => x(2),
				src(23) => x(1),
				src(24) => x(0),
				src(31 downto 25) => xin(31 downto 25),
	  			z => z(24)
				);
	mux_map25: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(25),
				src(1) => x(24),
				src(2) => x(23),
				src(3) => x(22),
				src(4) => x(21),
				src(5) => x(20),
				src(6) => x(19),
				src(7) => x(18),
				src(8) => x(17),
				src(9) => x(16),
				src(10) => x(15),
				src(11) => x(14),
				src(12) => x(13),
				src(13) => x(12),
				src(14) => x(11),
				src(15) => x(10),
				src(16) => x(9),
				src(17) => x(8),
				src(18) => x(7),
				src(19) => x(6),
				src(20) => x(5),
				src(21) => x(4),
				src(22) => x(3),
				src(23) => x(2),
				src(24) => x(1),
				src(25) => x(0),
				src(31 downto 26) => xin(31 downto 26),
	  			z => z(25)
				);
	mux_map26: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(26),
				src(1) => x(25),
				src(2) => x(24),
				src(3) => x(23),
				src(4) => x(22),
				src(5) => x(21),
				src(6) => x(20),
				src(7) => x(19),
				src(8) => x(18),
				src(9) => x(17),
				src(10) => x(16),
				src(11) => x(15),
				src(12) => x(14),
				src(13) => x(13),
				src(14) => x(12),
				src(15) => x(11),
				src(16) => x(10),
				src(17) => x(9),
				src(18) => x(8),
				src(19) => x(7),
				src(20) => x(6),
				src(21) => x(5),
				src(22) => x(4),
				src(23) => x(3),
				src(24) => x(2),
				src(25) => x(1),
				src(26) => x(0),
				src(31 downto 27) => xin(31 downto 27),
	  			z => z(26)
				);
	mux_map27: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(27),
				src(1) => x(26),
				src(2) => x(25),
				src(3) => x(24),
				src(4) => x(23),
				src(5) => x(22),
				src(6) => x(21),
				src(7) => x(20),
				src(8) => x(19),
				src(9) => x(18),
				src(10) => x(17),
				src(11) => x(16),
				src(12) => x(15),
				src(13) => x(14),
				src(14) => x(13),
				src(15) => x(12),
				src(16) => x(11),
				src(17) => x(10),
				src(18) => x(9),
				src(19) => x(8),
				src(20) => x(7),
				src(21) => x(6),
				src(22) => x(5),
				src(23) => x(4),
				src(24) => x(3),
				src(25) => x(2),
				src(26) => x(1),
				src(27) => x(0),
				src(31 downto 28) => xin(31 downto 28),
	  			z => z(27)
				);
	mux_map28: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(28),
				src(1) => x(27),
				src(2) => x(26),
				src(3) => x(25),
				src(4) => x(24),
				src(5) => x(23),
				src(6) => x(22),
				src(7) => x(21),
				src(8) => x(20),
				src(9) => x(19),
				src(10) => x(18),
				src(11) => x(17),
				src(12) => x(16),
				src(13) => x(15),
				src(14) => x(14),
				src(15) => x(13),
				src(16) => x(12),
				src(17) => x(11),
				src(18) => x(10),
				src(19) => x(9),
				src(20) => x(8),
				src(21) => x(7),
				src(22) => x(6),
				src(23) => x(5),
				src(24) => x(4),
				src(25) => x(3),
				src(26) => x(2),
				src(27) => x(1),
				src(28) => x(0),
				src(31 downto 29) => xin(31 downto 29),
	  			z => z(28)
				);
	mux_map29: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(29),
				src(1) => x(28),
				src(2) => x(27),
				src(3) => x(26),
				src(4) => x(25),
				src(5) => x(24),
				src(6) => x(23),
				src(7) => x(22),
				src(8) => x(21),
				src(9) => x(20),
				src(10) => x(19),
				src(11) => x(18),
				src(12) => x(17),
				src(13) => x(16),
				src(14) => x(15),
				src(15) => x(14),
				src(16) => x(13),
				src(17) => x(12),
				src(18) => x(11),
				src(19) => x(10),
				src(20) => x(9),
				src(21) => x(8),
				src(22) => x(7),
				src(23) => x(6),
				src(24) => x(5),
				src(25) => x(4),
				src(26) => x(3),
				src(27) => x(2),
				src(28) => x(1),
				src(29) => x(0),
				src(31 downto 30) => xin(31 downto 30),
	  			z => z(29)
				);
	mux_map30: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(30),
				src(1) => x(29),
				src(2) => x(28),
				src(3) => x(27),
				src(4) => x(26),
				src(5) => x(25),
				src(6) => x(24),
				src(7) => x(23),
				src(8) => x(22),
				src(9) => x(21),
				src(10) => x(20),
				src(11) => x(19),
				src(12) => x(18),
				src(13) => x(17),
				src(14) => x(16),
				src(15) => x(15),
				src(16) => x(14),
				src(17) => x(13),
				src(18) => x(12),
				src(19) => x(11),
				src(20) => x(10),
				src(21) => x(9),
				src(22) => x(8),
				src(23) => x(7),
				src(24) => x(6),
				src(25) => x(5),
				src(26) => x(4),
				src(27) => x(3),
				src(28) => x(2),
				src(29) => x(1),
				src(30) => x(0),
				src(31) => xin(31),
	  			z => z(30)
				);
	mux_map31: mux_32to1 port map (
	 		 	sel => shift (4 downto 0),
	  			src(0) => x(31),
				src(1) => x(30),
				src(2) => x(29),
				src(3) => x(28),
				src(4) => x(27),
				src(5) => x(26),
				src(6) => x(25),
				src(7) => x(24),
				src(8) => x(23),
				src(9) => x(22),
				src(10) => x(21),
				src(11) => x(20),
				src(12) => x(19),
				src(13) => x(18),
				src(14) => x(17),
				src(15) => x(16),
				src(16) => x(15),
				src(17) => x(14),
				src(18) => x(13),
				src(19) => x(12),
				src(20) => x(11),
				src(21) => x(10),
				src(22) => x(9),
				src(23) => x(8),
				src(24) => x(7),
				src(25) => x(6),
				src(26) => x(5),
				src(27) => x(4),
				src(28) => x(3),
				src(29) => x(2),
				src(30) => x(1),
				src(31) => x(0),
	  			z => z(31)
				);
end architecture structural;
